* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt custom_dff CLK D VGND VNB VPB VPWR Q
M0 a_891_413# a_193_47# a_975_413# VPB pfet_01v8_hvt w=0.42u l=0.15u
M1 a_1059_315# a_891_413# VGND VNB nfet_01v8 w=0.65u l=0.15u
M2 a_466_413# a_27_47# a_561_413# VPB pfet_01v8_hvt w=0.42u l=0.15u
M3 a_634_159# a_27_47# a_891_413# VPB pfet_01v8_hvt w=0.42u l=0.15u
M4 a_381_47# a_193_47# a_466_413# VPB pfet_01v8_hvt w=0.42u l=0.15u
M5 VPWR D a_381_47# VPB pfet_01v8_hvt w=0.42u l=0.15u
M6 VPWR a_466_413# a_634_159# VPB pfet_01v8_hvt w=0.75u l=0.15u
M7 VGND a_466_413# a_634_159# VNB nfet_01v8 w=0.64u l=0.15u
M8 a_1017_47# a_1059_315# VGND VNB nfet_01v8 w=0.42u l=0.15u
M9 a_1059_315# a_891_413# VPWR VPB pfet_01v8_hvt w=1u l=0.15u
M10 a_561_413# a_634_159# VPWR VPB pfet_01v8_hvt w=0.42u l=0.15u
M11 VPWR a_1059_315# Q VPB pfet_01v8_hvt w=1u l=0.15u
M12 a_891_413# a_27_47# a_1017_47# VNB nfet_01v8 w=0.36u l=0.15u
M13 a_634_159# a_193_47# a_891_413# VNB nfet_01v8 w=0.36u l=0.15u
M14 a_592_47# a_634_159# VGND VNB nfet_01v8 w=0.42u l=0.15u
M15 a_466_413# a_193_47# a_592_47# VNB nfet_01v8 w=0.36u l=0.15u
M16 VGND a_27_47# a_193_47# VNB nfet_01v8 w=0.42u l=0.15u
M17 a_381_47# a_27_47# a_466_413# VNB nfet_01v8 w=0.36u l=0.15u
M18 a_27_47# CLK VGND VNB nfet_01v8 w=0.42u l=0.15u
M19 a_27_47# CLK VPWR VPB pfet_01v8_hvt w=0.64u l=0.15u
M20 VPWR a_27_47# a_193_47# VPB pfet_01v8_hvt w=0.64u l=0.15u
M21 VGND D a_381_47# VNB nfet_01v8 w=0.42u l=0.15u
M22 a_975_413# a_1059_315# VPWR VPB pfet_01v8_hvt w=0.42u l=0.15u
M23 VGND a_1059_315# Q VNB nfet_01v8 w=0.65u l=0.15u
.ends
